module execute();



endmodule